module tb_full_subtractor();
    logic A, B, Bin;
    logic Diff, Bout;

    full_subtractor uut(A, B, Bin, Diff, Bout);

    initial begin
        A = 0; B = 0; Bin = 0; #10;
        A = 0; B = 0; Bin = 1; #10;
        A = 0; B = 1; Bin = 0; #10;
        A = 0; B = 1; Bin = 1; #10;
        A = 1; B = 0; Bin = 0; #10;
        A = 1; B = 0; Bin = 1; #10;
        A = 1; B = 1; Bin = 0; #10;
        A = 1; B = 1; Bin = 1; #10;
    end
endmodule
