module tb_johnson_counter;
    logic clock, reset;
    logic [3:0] q;

    johnson_counter dut (clock, reset, q);

    always #5 clock = ~clock;

    initial begin
        clock = 0; reset = 1;
        #10 reset = 0;
        #100 reset = 1;
        #10 reset = 0;
        #100 $stop;
    end
endmodule
